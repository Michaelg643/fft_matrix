type lut is array (natural range 0 to 510) of std_logic_vector(15 downto 0);
constant window_coe : lut := (
"0000000000001100",
"0000000000001110",
"0000000000010001",
"0000000000010101",
"0000000000011001",
"0000000000011101",
"0000000000100001",
"0000000000100110",
"0000000000101011",
"0000000000110001",
"0000000000110111",
"0000000000111110",
"0000000001000101",
"0000000001001101",
"0000000001010110",
"0000000001011111",
"0000000001101001",
"0000000001110011",
"0000000001111110",
"0000000010001010",
"0000000010010111",
"0000000010100100",
"0000000010110011",
"0000000011000010",
"0000000011010010",
"0000000011100011",
"0000000011110101",
"0000000100001001",
"0000000100011101",
"0000000100110010",
"0000000101001001",
"0000000101100001",
"0000000101111010",
"0000000110010100",
"0000000110110000",
"0000000111001101",
"0000000111101100",
"0000001000001100",
"0000001000101110",
"0000001001010001",
"0000001001110110",
"0000001010011100",
"0000001011000101",
"0000001011101111",
"0000001100011011",
"0000001101001001",
"0000001101111001",
"0000001110101011",
"0000001111011111",
"0000010000010101",
"0000010001001101",
"0000010010001000",
"0000010011000101",
"0000010100000100",
"0000010101000110",
"0000010110001010",
"0000010111010001",
"0000011000011010",
"0000011001100110",
"0000011010110101",
"0000011100000111",
"0000011101011011",
"0000011110110011",
"0000100000001101",
"0000100001101010",
"0000100011001011",
"0000100100101111",
"0000100110010101",
"0000101000000000",
"0000101001101101",
"0000101011011110",
"0000101101010011",
"0000101111001011",
"0000110001000110",
"0000110011000110",
"0000110101001001",
"0000110111001111",
"0000111001011010",
"0000111011101000",
"0000111101111011",
"0001000000010001",
"0001000010101100",
"0001000101001010",
"0001000111101101",
"0001001010010100",
"0001001101000000",
"0001001111101111",
"0001010010100011",
"0001010101011100",
"0001011000011001",
"0001011011011010",
"0001011110100000",
"0001100001101011",
"0001100100111010",
"0001101000001110",
"0001101011100111",
"0001101111000100",
"0001110010100111",
"0001110110001110",
"0001111001111010",
"0001111101101011",
"0010000001100001",
"0010000101011100",
"0010001001011011",
"0010001101100000",
"0010010001101010",
"0010010101111001",
"0010011010001101",
"0010011110100111",
"0010100011000101",
"0010100111101000",
"0010101100010001",
"0010110000111111",
"0010110101110001",
"0010111010101001",
"0010111111100110",
"0011000100101001",
"0011001001110000",
"0011001110111100",
"0011010100001110",
"0011011001100101",
"0011011111000000",
"0011100100100001",
"0011101010000111",
"0011101111110010",
"0011110101100010",
"0011111011010111",
"0100000001010000",
"0100000111001111",
"0100001101010010",
"0100010011011010",
"0100011001100111",
"0100011111111001",
"0100100110001111",
"0100101100101010",
"0100110011001010",
"0100111001101110",
"0101000000010110",
"0101000111000010",
"0101001101110011",
"0101010100101001",
"0101011011100010",
"0101100010011111",
"0101101001100000",
"0101110000100110",
"0101110111101110",
"0101111110111011",
"0110000110001011",
"0110001101011111",
"0110010100110110",
"0110011100010001",
"0110100011101110",
"0110101011001111",
"0110110010110011",
"0110111010011010",
"0111000010000011",
"0111001001101111",
"0111010001011110",
"0111011001001111",
"0111100001000010",
"0111101000110111",
"0111110000101110",
"0111111000101000",
"1000000000100011",
"1000001000011111",
"1000010000011101",
"1000011000011100",
"1000100000011101",
"1000101000011110",
"1000110000100000",
"1000111000100011",
"1001000000100111",
"1001001000101011",
"1001010000101111",
"1001011000110011",
"1001100000110111",
"1001101000111011",
"1001110000111111",
"1001111001000010",
"1010000001000100",
"1010001001000101",
"1010010001000101",
"1010011001000100",
"1010100001000010",
"1010101000111110",
"1010110000111000",
"1010111000110000",
"1011000000100110",
"1011001000011010",
"1011010000001100",
"1011010111111011",
"1011011111100111",
"1011100111001111",
"1011101110110101",
"1011110110011000",
"1011111101110111",
"1100000101010010",
"1100001100101010",
"1100010011111101",
"1100011011001100",
"1100100010010111",
"1100101001011101",
"1100110000011111",
"1100110111011011",
"1100111110010011",
"1101000101000101",
"1101001011110010",
"1101010010011010",
"1101011000111011",
"1101011111010111",
"1101100101101101",
"1101101011111100",
"1101110010000101",
"1101111000001000",
"1101111110000100",
"1110000011111001",
"1110001001100111",
"1110001111001110",
"1110010100101110",
"1110011010000110",
"1110011111010111",
"1110100100100000",
"1110101001100001",
"1110101110011011",
"1110110011001100",
"1110110111110101",
"1110111100010110",
"1111000000101110",
"1111000100111110",
"1111001001000101",
"1111001101000011",
"1111010000111000",
"1111010100100101",
"1111011000001000",
"1111011011100010",
"1111011110110011",
"1111100001111010",
"1111100100111000",
"1111100111101101",
"1111101010011000",
"1111101100111001",
"1111101111010000",
"1111110001011110",
"1111110011100010",
"1111110101011100",
"1111110111001100",
"1111111000110001",
"1111111010001101",
"1111111011011111",
"1111111100100111",
"1111111101100100",
"1111111110010111",
"1111111111000000",
"1111111111011111",
"1111111111110011",
"1111111111111110",
"1111111111111110",
"1111111111110011",
"1111111111011111",
"1111111111000000",
"1111111110010111",
"1111111101100100",
"1111111100100111",
"1111111011011111",
"1111111010001101",
"1111111000110001",
"1111110111001100",
"1111110101011100",
"1111110011100010",
"1111110001011110",
"1111101111010000",
"1111101100111001",
"1111101010011000",
"1111100111101101",
"1111100100111000",
"1111100001111010",
"1111011110110011",
"1111011011100010",
"1111011000001000",
"1111010100100101",
"1111010000111000",
"1111001101000011",
"1111001001000101",
"1111000100111110",
"1111000000101110",
"1110111100010110",
"1110110111110101",
"1110110011001100",
"1110101110011011",
"1110101001100001",
"1110100100100000",
"1110011111010111",
"1110011010000110",
"1110010100101110",
"1110001111001110",
"1110001001100111",
"1110000011111001",
"1101111110000100",
"1101111000001000",
"1101110010000101",
"1101101011111100",
"1101100101101101",
"1101011111010111",
"1101011000111011",
"1101010010011010",
"1101001011110010",
"1101000101000101",
"1100111110010011",
"1100110111011011",
"1100110000011111",
"1100101001011101",
"1100100010010111",
"1100011011001100",
"1100010011111101",
"1100001100101010",
"1100000101010010",
"1011111101110111",
"1011110110011000",
"1011101110110101",
"1011100111001111",
"1011011111100111",
"1011010111111011",
"1011010000001100",
"1011001000011010",
"1011000000100110",
"1010111000110000",
"1010110000111000",
"1010101000111110",
"1010100001000010",
"1010011001000100",
"1010010001000101",
"1010001001000101",
"1010000001000100",
"1001111001000010",
"1001110000111111",
"1001101000111011",
"1001100000110111",
"1001011000110011",
"1001010000101111",
"1001001000101011",
"1001000000100111",
"1000111000100011",
"1000110000100000",
"1000101000011110",
"1000100000011101",
"1000011000011100",
"1000010000011101",
"1000001000011111",
"1000000000100011",
"0111111000101000",
"0111110000101110",
"0111101000110111",
"0111100001000010",
"0111011001001111",
"0111010001011110",
"0111001001101111",
"0111000010000011",
"0110111010011010",
"0110110010110011",
"0110101011001111",
"0110100011101110",
"0110011100010001",
"0110010100110110",
"0110001101011111",
"0110000110001011",
"0101111110111011",
"0101110111101110",
"0101110000100110",
"0101101001100000",
"0101100010011111",
"0101011011100010",
"0101010100101001",
"0101001101110011",
"0101000111000010",
"0101000000010110",
"0100111001101110",
"0100110011001010",
"0100101100101010",
"0100100110001111",
"0100011111111001",
"0100011001100111",
"0100010011011010",
"0100001101010010",
"0100000111001111",
"0100000001010000",
"0011111011010111",
"0011110101100010",
"0011101111110010",
"0011101010000111",
"0011100100100001",
"0011011111000000",
"0011011001100101",
"0011010100001110",
"0011001110111100",
"0011001001110000",
"0011000100101001",
"0010111111100110",
"0010111010101001",
"0010110101110001",
"0010110000111111",
"0010101100010001",
"0010100111101000",
"0010100011000101",
"0010011110100111",
"0010011010001101",
"0010010101111001",
"0010010001101010",
"0010001101100000",
"0010001001011011",
"0010000101011100",
"0010000001100001",
"0001111101101011",
"0001111001111010",
"0001110110001110",
"0001110010100111",
"0001101111000100",
"0001101011100111",
"0001101000001110",
"0001100100111010",
"0001100001101011",
"0001011110100000",
"0001011011011010",
"0001011000011001",
"0001010101011100",
"0001010010100011",
"0001001111101111",
"0001001101000000",
"0001001010010100",
"0001000111101101",
"0001000101001010",
"0001000010101100",
"0001000000010001",
"0000111101111011",
"0000111011101000",
"0000111001011010",
"0000110111001111",
"0000110101001001",
"0000110011000110",
"0000110001000110",
"0000101111001011",
"0000101101010011",
"0000101011011110",
"0000101001101101",
"0000101000000000",
"0000100110010101",
"0000100100101111",
"0000100011001011",
"0000100001101010",
"0000100000001101",
"0000011110110011",
"0000011101011011",
"0000011100000111",
"0000011010110101",
"0000011001100110",
"0000011000011010",
"0000010111010001",
"0000010110001010",
"0000010101000110",
"0000010100000100",
"0000010011000101",
"0000010010001000",
"0000010001001101",
"0000010000010101",
"0000001111011111",
"0000001110101011",
"0000001101111001",
"0000001101001001",
"0000001100011011",
"0000001011101111",
"0000001011000101",
"0000001010011100",
"0000001001110110",
"0000001001010001",
"0000001000101110",
"0000001000001100",
"0000000111101100",
"0000000111001101",
"0000000110110000",
"0000000110010100",
"0000000101111010",
"0000000101100001",
"0000000101001001",
"0000000100110010",
"0000000100011101",
"0000000100001001",
"0000000011110101",
"0000000011100011",
"0000000011010010",
"0000000011000010",
"0000000010110011",
"0000000010100100",
"0000000010010111",
"0000000010001010",
"0000000001111110",
"0000000001110011",
"0000000001101001",
"0000000001011111",
"0000000001010110",
"0000000001001101",
"0000000001000101",
"0000000000111110",
"0000000000110111",
"0000000000110001",
"0000000000101011",
"0000000000100110",
"0000000000100001",
"0000000000011101",
"0000000000011001",
"0000000000010101",
"0000000000010001",
"0000000000001110");
