type lut is array (natural range 0 to 254) of std_logic_vector(15 downto 0);
constant window_coe : lut := (
"0000000000001100",
"0000000000010001",
"0000000000011001",
"0000000000100001",
"0000000000101100",
"0000000000111000",
"0000000001000110",
"0000000001010111",
"0000000001101010",
"0000000001111111",
"0000000010011000",
"0000000010110101",
"0000000011010101",
"0000000011111000",
"0000000100100000",
"0000000101001101",
"0000000101111111",
"0000000110110110",
"0000000111110011",
"0000001000110101",
"0000001001111111",
"0000001011001111",
"0000001100100111",
"0000001110000110",
"0000001111101110",
"0000010001011110",
"0000010011011000",
"0000010101011011",
"0000010111101001",
"0000011010000001",
"0000011100100100",
"0000011111010011",
"0000100010001110",
"0000100101010110",
"0000101000101011",
"0000101100001110",
"0000101111111111",
"0000110011111110",
"0000111000001101",
"0000111100101011",
"0001000001011010",
"0001000110011001",
"0001001011101001",
"0001010001001010",
"0001010110111101",
"0001011101000011",
"0001100011011011",
"0001101010000110",
"0001110001000100",
"0001111000010110",
"0001111111111011",
"0010000111110101",
"0010010000000011",
"0010011000100110",
"0010100001011101",
"0010101010101000",
"0010110100001001",
"0010111101111110",
"0011001000001000",
"0011010010100111",
"0011011101011011",
"0011101000100011",
"0011110011111111",
"0011111111101111",
"0100001011110011",
"0100011000001011",
"0100100100110101",
"0100110001110011",
"0100111111000010",
"0101001100100011",
"0101011010010101",
"0101101000011000",
"0101110110101010",
"0110000101001011",
"0110010011111011",
"0110100010111000",
"0110110010000001",
"0111000001010111",
"0111010000110111",
"0111100000100000",
"0111110000010011",
"1000000000001101",
"1000010000001101",
"1000100000010011",
"1000110000011100",
"1001000000101001",
"1001010000110111",
"1001100001000110",
"1001110001010011",
"1010000001011110",
"1010010001100110",
"1010100001101000",
"1010110001100100",
"1011000001011000",
"1011010001000010",
"1011100000100010",
"1011101111110110",
"1011111110111100",
"1100001101110011",
"1100011100011010",
"1100101010101111",
"1100111000110001",
"1101000110011110",
"1101010011110101",
"1101100000110100",
"1101101101011011",
"1101111001101000",
"1110000101011010",
"1110010000110000",
"1110011011101000",
"1110100110000001",
"1110101111111010",
"1110111001010011",
"1111000010001010",
"1111001010011110",
"1111010010001110",
"1111011001011010",
"1111100000000000",
"1111100110000000",
"1111101011011010",
"1111110000001101",
"1111110100010111",
"1111110111111010",
"1111111010110100",
"1111111101000100",
"1111111110101100",
"1111111111101010",
"1111111111111111",
"1111111111101010",
"1111111110101100",
"1111111101000100",
"1111111010110100",
"1111110111111010",
"1111110100010111",
"1111110000001101",
"1111101011011010",
"1111100110000000",
"1111100000000000",
"1111011001011010",
"1111010010001110",
"1111001010011110",
"1111000010001010",
"1110111001010011",
"1110101111111010",
"1110100110000001",
"1110011011101000",
"1110010000110000",
"1110000101011010",
"1101111001101000",
"1101101101011011",
"1101100000110100",
"1101010011110101",
"1101000110011110",
"1100111000110001",
"1100101010101111",
"1100011100011010",
"1100001101110011",
"1011111110111100",
"1011101111110110",
"1011100000100010",
"1011010001000010",
"1011000001011000",
"1010110001100100",
"1010100001101000",
"1010010001100110",
"1010000001011110",
"1001110001010011",
"1001100001000110",
"1001010000110111",
"1001000000101001",
"1000110000011100",
"1000100000010011",
"1000010000001101",
"1000000000001101",
"0111110000010011",
"0111100000100000",
"0111010000110111",
"0111000001010111",
"0110110010000001",
"0110100010111000",
"0110010011111011",
"0110000101001011",
"0101110110101010",
"0101101000011000",
"0101011010010101",
"0101001100100011",
"0100111111000010",
"0100110001110011",
"0100100100110101",
"0100011000001011",
"0100001011110011",
"0011111111101111",
"0011110011111111",
"0011101000100011",
"0011011101011011",
"0011010010100111",
"0011001000001000",
"0010111101111110",
"0010110100001001",
"0010101010101000",
"0010100001011101",
"0010011000100110",
"0010010000000011",
"0010000111110101",
"0001111111111011",
"0001111000010110",
"0001110001000100",
"0001101010000110",
"0001100011011011",
"0001011101000011",
"0001010110111101",
"0001010001001010",
"0001001011101001",
"0001000110011001",
"0001000001011010",
"0000111100101011",
"0000111000001101",
"0000110011111110",
"0000101111111111",
"0000101100001110",
"0000101000101011",
"0000100101010110",
"0000100010001110",
"0000011111010011",
"0000011100100100",
"0000011010000001",
"0000010111101001",
"0000010101011011",
"0000010011011000",
"0000010001011110",
"0000001111101110",
"0000001110000110",
"0000001100100111",
"0000001011001111",
"0000001001111111",
"0000001000110101",
"0000000111110011",
"0000000110110110",
"0000000101111111",
"0000000101001101",
"0000000100100000",
"0000000011111000",
"0000000011010101",
"0000000010110101",
"0000000010011000",
"0000000001111111",
"0000000001101010",
"0000000001010111",
"0000000001000110",
"0000000000111000",
"0000000000101100",
"0000000000100001",
"0000000000011001",
"0000000000010001",
"0000000000001100");
