type lut is array (natural range 0 to 254) of std_logic_vector(15 downto 0);
constant window_coe : lut := (
"0000000000001100",
"0000000000010001",
"0000000000011001",
"0000000000100001",
"0000000000101011",
"0000000000110111",
"0000000001000110",
"0000000001010110",
"0000000001101001",
"0000000001111111",
"0000000010010111",
"0000000010110011",
"0000000011010011",
"0000000011110110",
"0000000100011110",
"0000000101001010",
"0000000101111100",
"0000000110110010",
"0000000111101110",
"0000001000110000",
"0000001001111001",
"0000001011001000",
"0000001100011111",
"0000001101111101",
"0000001111100100",
"0000010001010011",
"0000010011001011",
"0000010101001101",
"0000010111011001",
"0000011001101111",
"0000011100010000",
"0000011110111101",
"0000100001110110",
"0000100100111100",
"0000101000001110",
"0000101011101110",
"0000101111011100",
"0000110011011000",
"0000110111100100",
"0000111011111111",
"0001000000101001",
"0001000101100100",
"0001001010110000",
"0001010000001101",
"0001010101111100",
"0001011011111101",
"0001100010010000",
"0001101000110110",
"0001101111101110",
"0001110110111011",
"0001111110011011",
"0010000110001110",
"0010001110010110",
"0010010110110010",
"0010011111100011",
"0010101000101000",
"0010110010000010",
"0010111011110000",
"0011000101110011",
"0011010000001010",
"0011011010110110",
"0011100101110110",
"0011110001001011",
"0011111100110011",
"0100001000110000",
"0100010100111111",
"0100100001100010",
"0100101110010111",
"0100111011011110",
"0101001000110111",
"0101010110100001",
"0101100100011100",
"0101110010100110",
"0110000001000000",
"0110001111101000",
"0110011110011101",
"0110101101011111",
"0110111100101101",
"0111001100000110",
"0111011011101001",
"0111101011010101",
"0111111011001000",
"1000001011000011",
"1000011011000011",
"1000101011000111",
"1000111011001111",
"1001001011011001",
"1001011011100011",
"1001101011101101",
"1001111011110101",
"1010001011111010",
"1010011011111010",
"1010101011110101",
"1010111011101000",
"1011001011010010",
"1011011010110010",
"1011101010000111",
"1011111001001110",
"1100001000001000",
"1100010110110001",
"1100100101001010",
"1100110011001111",
"1101000001000001",
"1101001110011110",
"1101011011100100",
"1101101000010010",
"1101110100100111",
"1110000000100001",
"1110001100000000",
"1110010111000010",
"1110100001100110",
"1110101011101011",
"1110110101001111",
"1110111110010011",
"1111000110110100",
"1111001110110011",
"1111010110001101",
"1111011101000011",
"1111100011010011",
"1111101000111110",
"1111101110000001",
"1111110010011110",
"1111110110010010",
"1111111001011111",
"1111111100000011",
"1111111101111110",
"1111111111010001",
"1111111111111010",
"1111111111111010",
"1111111111010001",
"1111111101111110",
"1111111100000011",
"1111111001011111",
"1111110110010010",
"1111110010011110",
"1111101110000001",
"1111101000111110",
"1111100011010011",
"1111011101000011",
"1111010110001101",
"1111001110110011",
"1111000110110100",
"1110111110010011",
"1110110101001111",
"1110101011101011",
"1110100001100110",
"1110010111000010",
"1110001100000000",
"1110000000100001",
"1101110100100111",
"1101101000010010",
"1101011011100100",
"1101001110011110",
"1101000001000001",
"1100110011001111",
"1100100101001010",
"1100010110110001",
"1100001000001000",
"1011111001001110",
"1011101010000111",
"1011011010110010",
"1011001011010010",
"1010111011101000",
"1010101011110101",
"1010011011111010",
"1010001011111010",
"1001111011110101",
"1001101011101101",
"1001011011100011",
"1001001011011001",
"1000111011001111",
"1000101011000111",
"1000011011000011",
"1000001011000011",
"0111111011001000",
"0111101011010101",
"0111011011101001",
"0111001100000110",
"0110111100101101",
"0110101101011111",
"0110011110011101",
"0110001111101000",
"0110000001000000",
"0101110010100110",
"0101100100011100",
"0101010110100001",
"0101001000110111",
"0100111011011110",
"0100101110010111",
"0100100001100010",
"0100010100111111",
"0100001000110000",
"0011111100110011",
"0011110001001011",
"0011100101110110",
"0011011010110110",
"0011010000001010",
"0011000101110011",
"0010111011110000",
"0010110010000010",
"0010101000101000",
"0010011111100011",
"0010010110110010",
"0010001110010110",
"0010000110001110",
"0001111110011011",
"0001110110111011",
"0001101111101110",
"0001101000110110",
"0001100010010000",
"0001011011111101",
"0001010101111100",
"0001010000001101",
"0001001010110000",
"0001000101100100",
"0001000000101001",
"0000111011111111",
"0000110111100100",
"0000110011011000",
"0000101111011100",
"0000101011101110",
"0000101000001110",
"0000100100111100",
"0000100001110110",
"0000011110111101",
"0000011100010000",
"0000011001101111",
"0000010111011001",
"0000010101001101",
"0000010011001011",
"0000010001010011",
"0000001111100100",
"0000001101111101",
"0000001100011111",
"0000001011001000",
"0000001001111001",
"0000001000110000",
"0000000111101110",
"0000000110110010",
"0000000101111100",
"0000000101001010",
"0000000100011110",
"0000000011110110",
"0000000011010011",
"0000000010110011",
"0000000010010111",
"0000000001111111",
"0000000001101001",
"0000000001010110",
"0000000001000110",
"0000000000110111",
"0000000000101011",
"0000000000100001",
"0000000000011001",
"0000000000010001");
